library verilog;
use verilog.vl_types.all;
entity BANCOdeREGISTRADORES32bits_vlg_vec_tst is
end BANCOdeREGISTRADORES32bits_vlg_vec_tst;
