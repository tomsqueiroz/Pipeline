library verilog;
use verilog.vl_types.all;
entity TESTE_vlg_vec_tst is
end TESTE_vlg_vec_tst;
